library verilog;
use verilog.vl_types.all;
entity testing_reg_tb is
end testing_reg_tb;
