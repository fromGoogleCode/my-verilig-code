library verilog;
use verilog.vl_types.all;
entity nand_write_tb is
end nand_write_tb;
