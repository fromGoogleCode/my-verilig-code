library verilog;
use verilog.vl_types.all;
entity my_toggle_tb is
end my_toggle_tb;
