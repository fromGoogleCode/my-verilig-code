library verilog;
use verilog.vl_types.all;
entity my_pll_tb is
end my_pll_tb;
