library verilog;
use verilog.vl_types.all;
entity readID_tb is
end readID_tb;
